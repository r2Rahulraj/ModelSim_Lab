module ha_st(s,c,a,b);
input a,b;
output c,s;

and a1(c,a,b);
or o1(s,a,b);

endmodule